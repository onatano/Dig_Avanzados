library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.numeric_std.all;

entity Deco is
    port (
        stage : in std_logic_vector(2 downto 0);
        clear,enable,store : out std_logic
	);
end entity;

architecture Beh of Deco is

    begin

       
    
end Beh;